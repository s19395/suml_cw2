���,      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.0.1�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�auto�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�objawy��wiek��choroby��wzrost�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��h2�f8�����R�(KhHNNNJ����J����K t�b�C              �?�t�bhLh&�scalar���hGC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hK�
node_count�K�nodes�h(h+K ��h-��R�(KK��h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hxhGK ��hyhGK��hzhGK��h{hXK��h|hXK ��h}hGK(��h~hXK0��uK8KKt�b�B                              @|��?���?"             K@                           @ܷ��?��?             =@������������������������       �                     :@������������������������       �                     @������������������������       �                     9@�t�b�values�h(h+K ��h-��R�(KKKK��hX�CP      :@      <@      :@      @      :@                      @              9@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�BH                              @      �?$             K@                            @     ��?             @@������������������������       �                     5@                          �g@�eP*L��?	             &@                          �E@����X�?             @                          �:@      �?             @������������������������       �                     �?                           �?�q�q�?             @	       
                   �@@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     6@�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      ;@      ;@      ;@      @      5@              @      @       @      @       @       @              �?       @      �?      �?      �?      �?                      �?      �?                      @      @                      6@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                              @      �?!             K@������������������������       �                     7@       
                   �h@��� ��?             ?@                          �g@ ��WV�?             :@������������������������       �        
             6@       	                    h@      �?             @                            @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                            @���Q��?             @������������������������       �                     @������������������������       �                      @�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      ;@      ;@      7@              @      ;@      �?      9@              6@      �?      @      �?      �?      �?                      �?               @      @       @      @                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                              @|��?���?!             K@                            @��S�ۿ?             >@������������������������       �                     8@                         �f@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     8@�t�bh�h(h+K ��h-��R�(KKKK��hX�Cp      <@      :@      <@       @      8@              @       @               @      @                      8@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoK	hph(h+K ��h-��R�(KK	��hw�B�                              @���3L�?'             K@������������������������       �                     4@                            @l��\��?             A@                           @      �?              @                         ��e@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     :@�t�bh�h(h+K ��h-��R�(KK	KK��hX�C�      7@      ?@      4@              @      ?@      @      @      @       @               @      @                      @              :@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoK	hph(h+K ��h-��R�(KK	��hw�B�                            �d@�q�q�?#             K@������������������������       �                     @                           �?�t����?!            �I@                            @      �?             8@������������������������       �                     ,@                         y�E@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     ;@�t�bh�h(h+K ��h-��R�(KK	KK��hX�C�      2@      B@      @              .@      B@      .@      "@      ,@              �?      "@              "@      �?                      ;@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoK	hph(h+K ��h-��R�(KK	��hw�B�                            @E@�5��?!             K@                            @և���X�?             5@������������������������       �                     "@������������������������       �                     (@                            @:ɨ��?            �@@������������������������       �                     6@                           �?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KK	KK��hX�C�      @@      6@      "@      (@      "@                      (@      7@      $@      6@              �?      $@      �?                      $@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoK	hph(h+K ��h-��R�(KK	��hw�B�                              @�5��?$             K@������������������������       �                     4@                           @�IєX�?             A@                            @�����H�?             2@                           f@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �        	             ,@������������������������       �                     0@�t�bh�h(h+K ��h-��R�(KK	KK��hX�C�      6@      @@      4@               @      @@       @      0@       @       @               @       @                      ,@              0@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�Bh                            �f@b�2�tk�?$             K@                            @D�n�3�?             3@������������������������       �                     &@������������������������       �                      @                            @����X�?            �A@������������������������       �                     @       
                     @\-��p�?             =@       	                   �E@���Q��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     3@�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      5@     �@@      &@       @      &@                       @      $@      9@      @              @      9@      @      @      @                      @              3@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                              @�q�q�?             K@������������������������       �                     (@                           @؇���X�?             E@                            @�θ�?             :@                           f@      �?              @������������������������       �                     �?       
                   �g@؇���X�?             @       	                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �        	             2@������������������������       �                     0@�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      2@      B@      (@              @      B@      @      4@      @       @              �?      @      �?       @      �?              �?       @              @                      2@              0@�t�bubhhubehhub.